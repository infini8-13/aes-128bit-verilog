module ALL_ENC_TEST;

wire DONE,DONE1,DONE2,DONE3;
reg RST,CLK;
/*
CIPHER_FEEDBACK_MODE_ENC M1(DONE,CLK,RST);
CIPHER_CHAINING_MODE_ENC M2(DONE1,CLK,RST);
OUTPUT_FEEDBACK_MODE_ENC M3(DONE2,CLK,RST);
INDEX_MODE_ENC M4(DONE3,CLK,RST);
*/

INDEX_MODE_DEC M5(DONE,CLK,RST);
OUTPUT_FEEDBACK_MODE_DEC M6(DONE1,CLK,RST);
CIPHER_CHAINING_MODE_DEC M7(DONE2,CLK,RST);
CIPHER_FEEDBACK_MODE_DEC M8(DONE3,CLK,RST);


initial begin CLK=1'b0; RST=1'b0; #200 RST=1'b1; end
always #5 CLK=~CLK;

endmodule
