module KEY_GENERATOR(RK,GENERATED,UK,GENERATE,RST,CLK);

output reg[0:767] RK;
output reg GENERATED;
input [0:63]UK;
input GENERATE,RST,CLK;

reg [0:55]K;

always @(negedge CLK or negedge RST) 
if(~RST) begin GENERATED <= 1'b0; RK<=768'b0; K<=56'b0; end 
else if({GENERATE,GENERATED} == 2'b10) begin

K[0]=UK[56]   ; K[1]=UK[48]  ; K[2]=UK[40]  ; K[3]=UK[32]  ; K[4]=UK[24]  ; K[5]=UK[16]  ; K[6]=UK[8]   ;
K[7]=UK[0]   ; K[8]=UK[57]  ; K[9]=UK[49]  ; K[10]=UK[41] ; K[11]=UK[33] ; K[12]=UK[25] ; K[13]=UK[17] ;
K[14]=UK[9]  ; K[15]=UK[1]  ; K[16]=UK[58] ; K[17]=UK[50] ; K[18]=UK[42] ; K[19]=UK[34] ; K[20]=UK[26] ;
K[21]=UK[18] ; K[22]=UK[10] ; K[23]=UK[2]  ; K[24]=UK[59] ; K[25]=UK[51] ; K[26]=UK[43] ; K[27]=UK[35] ;
K[28]=UK[62] ; K[29]=UK[54] ; K[30]=UK[46] ; K[31]=UK[38] ; K[32]=UK[30] ; K[33]=UK[22] ; K[34]=UK[14] ;
K[35]=UK[6]  ; K[36]=UK[61] ; K[37]=UK[53] ; K[38]=UK[45] ; K[39]=UK[37] ; K[40]=UK[29] ; K[41]=UK[21] ;
K[42]=UK[13] ; K[43]=UK[5]  ; K[44]=UK[60] ; K[45]=UK[52] ; K[46]=UK[44] ; K[47]=UK[36] ; K[48]=UK[28] ;
K[49]=UK[20] ; K[50]=UK[12] ; K[51]=UK[4]  ; K[52]=UK[27] ; K[53]=UK[19] ; K[54]=UK[11] ; K[55]=UK[3]   ; 


K = {K[1:27],K[0],K[29:55],K[28]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};

K = {K[1:27],K[0],K[29:55],K[28]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};

K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   

K = {K[1:27],K[0],K[29:55],K[28]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   
   
K = {K[2:27],K[0:1],K[30:55],K[28:29]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;
RK = {RK[48:767],RK[0:47]};   

K = {K[1:27],K[0],K[29:55],K[28]};
RK[720]=K[13] ; RK[721]=K[16] ; RK[722]=K[10] ; RK[723]=K[23] ; RK[724]=K[0]  ; RK[725]=K[4]  ; RK[726]=K[2]  ; RK[727]=K[27] ;
RK[728]=K[14] ; RK[729]=K[5]  ; RK[730]=K[20] ; RK[731]=K[9]  ; RK[732]=K[22] ; RK[733]=K[18] ; RK[734]=K[11] ; RK[735]=K[3]  ;
RK[736]=K[25] ; RK[737]=K[7]  ; RK[738]=K[15] ; RK[739]=K[6]  ; RK[740]=K[26] ; RK[741]=K[19] ; RK[742]=K[12] ; RK[743]=K[1]  ;
RK[744]=K[40] ; RK[745]=K[51] ; RK[746]=K[30] ; RK[747]=K[36] ; RK[748]=K[46] ; RK[749]=K[54] ; RK[750]=K[29] ; RK[751]=K[39] ;
RK[752]=K[50] ; RK[753]=K[44] ; RK[754]=K[32] ; RK[755]=K[47] ; RK[756]=K[43] ; RK[757]=K[48] ; RK[758]=K[38] ; RK[759]=K[55] ;
RK[760]=K[33] ; RK[761]=K[52] ; RK[762]=K[45] ; RK[763]=K[41] ; RK[764]=K[49] ; RK[765]=K[35] ; RK[766]=K[28] ; RK[767]=K[31] ;

GENERATED <= 1'b1;

end

endmodule
